--------------------------------------------------------------------------------
-- Processor test bench
--

library ieee;
use ieee.std_logic_1164.ALL;
use ieee.numeric_std.all;
 
library work;
use work.asserts.all;
 
entity processor_tb is
end processor_tb;
 
architecture behavior of processor_tb is
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    component processor port (
         clk               : in std_logic;
         reset             : in  std_logic;
         processor_enable  : in  std_logic;
         imem_address      : out  std_logic_vector(31 downto 0);
         imem_data_in      : in  std_logic_vector(31 downto 0);
         dmem_data_in      : in  std_logic_vector(31 downto 0);
         dmem_address      : out  std_logic_vector(31 downto 0);
         dmem_address_wr   : out  std_logic_vector(31 downto 0);
         dmem_data_out     : out  std_logic_vector(31 downto 0);
         dmem_write_enable : out  std_logic
        );
    end component;
    

   --Inputs
   signal clk : std_logic := '0';
   signal reset : std_logic := '0';
   signal processor_enable : std_logic := '0';
   signal imem_data_in : std_logic_vector(31 downto 0) := (others => '0');
   signal dmem_data_in : std_logic_vector(31 downto 0) := (others => '0');

 	--Outputs
   signal imem_address : std_logic_vector(31 downto 0);
   signal dmem_address : std_logic_vector(31 downto 0);
   signal dmem_address_wr : std_logic_vector(31 downto 0);
   signal dmem_data_out : std_logic_vector(31 downto 0);
   signal dmem_write_enable : std_logic;

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
begin
 
	-- Instantiate the Unit Under Test (UUT)
   uut: processor port map (
          clk => clk,
          reset => reset,
          processor_enable => processor_enable,
          imem_address => imem_address,
          imem_data_in => imem_data_in,
          dmem_data_in => dmem_data_in,
          dmem_address => dmem_address,
          dmem_address_wr => dmem_address_wr,
          dmem_data_out => dmem_data_out,
          dmem_write_enable => dmem_write_enable
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '1';
		wait for clk_period/2;
		clk <= '0';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
		-- hold reset state for 100 ns.
		wait for 100 ns;	
		reset <= '0';
		processor_enable <= '1';

		-- imem_data_in <= "00010000001000000000000000000001"; -- jump

		-- Load data memory 0 (Set intruction, wait for execute, assert dbus address and then wait for fetch)
		imem_data_in <= "10001100001000010000000000000010";
		dmem_data_in <= "00000000000000000000000000000010";
		wait for clk_period*2;
		assertEqual(dmem_address, "00000000000000000000000000000010","00000000000000000000000000000010");
		wait for clk_period;

		-- Branch if r0 and r1 are equal (They should not be, so we expect program counter to be 8 in next fetch
		imem_data_in <= "00010000001000000000000000000001";
		wait for clk_period*2;
		assertEqual(imem_address, "00000000000000000000000000000100","00000000000000000000000000000100");

		-- Branch if r1 and r1 are equal (The are, so we expect program counter to be 16 during next fetch)
		imem_data_in <= "00010000001000010000000000000001";
		wait for clk_period*2;
		wait for clk_period/2;
		assertEqual(imem_address, "00000000000000000000000000010000","00000000000000000000000000010000");

		-- Load upper immediate (32 << 16)
		imem_data_in <= "00111100000000100000000000100000";
		wait for clk_period/2;
		wait for clk_period;

		-- Write r2 to memory to validate previous instruction
		imem_data_in <= "10101100000000100000000000000000";
		wait for clk_period*3;
		assertEqual(dmem_data_out, "00000000001000000000000000000000", "00000000001000000000000000000000");


		wait;
   end process;

end;
